//Created by Peter Johnson
//pjohnson@g.hmc.edu
//Sep 16 2018
//Summary control 2 7-segment displays using a single 7-bit decoder and time multiplexing
module lab2_PJ(input logic clk,
					input logic [3:0] s0,
					input logic [3:0] s1,
					output logic [1:0] anode, //turns anodes on and off, anode 1 correspons to s1 and display 1
					output logic [7:0] led,
					output logic [6:0] seg);
	//Internal Logic variables
	logic [3:0] s; //currently selected input
	logic [31:0] q; // word with most significant bit to be toggled
	logic cycle; //either on the 0 half cycle or the 1 half cycle
	
	//Operation will occur at 60Hz
	//Will use a counter module defined below
	counter countLED(clk, q); 
	
	//Cycle will toggle at the same freq as the most significant bit
	//0 Cycle is when s is s0, and display 0 is lit, 1 cycle is when s is s1 and display 1 is lit
	assign cycle=q[31];
	
	//Multiplex based on what cycle we are on
	mux2 timeMux(s0,s1,cycle,s);
	
	//Turn on the anode depedning on which half cycle is the current one
	assign anode[1]= cycle; //when cycle=1 turn anode[1] on
	assign anode[0]= ~cycle; //opposite for anode[0]
	
	//Display the sum of two hexadecimal numbers on led[7:3]
	assign led[7:3]=s0+s1; //implies a full adder in hardware
	
	//7 Segment display logic
	//Encoding-	 seg 6543210
	// 				  abcdefg
	always_comb
		case(s)
		4'b0000:seg=7'b0000001; //0
		4'b0001:seg=7'b1001111; //1
		4'b0010:seg=7'b0010010; //2
		4'b0011:seg=7'b0000110; //3
		4'b0100:seg=7'b1001100; //4
		4'b0101:seg=7'b0100100; //5
		4'b0110:seg=7'b0100000; //6
		4'b0111:seg=7'b0001111; //7
		4'b1000:seg=7'b0000000; //8
		4'b1001:seg=7'b0001100; //9
		4'b1010:seg=7'b0001000; //A
		4'b1011:seg=7'b1100000; //b
		4'b1100:seg=7'b0110001; //C
		4'b1101:seg=7'b1000010; //d
		4'b1110:seg=7'b0110000; //E
		4'b1111:seg=7'b0111000; //F
		default:seg=7'b0110110; //Default is to display 3 horizontal lines which should never happen-can tell something is wrong
		endcase
		
		//Note that to turn on the LEDs we actually need to pass a 0 not a 1 so truth table looks inverted from what it normally is
	
endmodule

//Idiomatic counter code provided by Prof David Harris in Ch. 5 slides
//Modified by Peter Johnson September 16, 2018
//pjohnson@g.hmc.edu
//a divide by 2^N counter where the most significant bit toggles every 2^N cycles
//value of p(value incremented) selected so that toggling occurs at 60 Hz.
//Value is 60Hz about the edge of what is visible for the human eye
//fout=fclk*p/2^N
//fout=60 Hz, fclk=40MHz, N=32 bits so p=6442
module counter (input logic clk,
					 output logic [31:0] q);
 always_ff @ (posedge clk)
				q <= q+6442;
		
endmodule

//Idiomatic 2:1 multiplexer using conditional assignment
//Provided by David Harris-Digital Design and Computer Architecture
module mux2 (input logic[3:0] d0,d1,
				input logic 		s,
				output logic[3:0] y);
	// if s=1 y=d1, if s=0, y=d0
	assign y=s?d1:d0;
endmodule


