/////////////////////////////////////////////
// VGA.sv
// HMC E155 15 November 2018
// pjohnson@g.hmc.edu @tdubno@g.hmc.edu
// For MicroP's Final Project
// Implements VGA driver that takes in the message to be displayed through spi
// Msg component displays on one line, location component displays on another line
/////////////////////////////////////////////


/////////////////////////////////////////////
// VGA
// Top level module with SPI interface and VGA core
/////////////////////////////////////////////
module VGA(input  logic clk, 				//From 40 MHz oscillator
           input  logic sck, 				//From Pi
           input  logic sdi, 				//From Pi
			  output logic hsync, vsync,	//To VGA cable
			  output logic r,g,b); 			//To vga cable
    
	 //intermdiate logic	 
    logic [15:0] received;					
	 logic [7:0] char;
	 logic vgaclk,done,clkdone,msgEn;
    
	 //instantiate spi module
    vga_spi spi(sck,sdi,done,received);   
	 assign char = received[7:0];			//2nd half of short is the char to be displayed
	 assign msgEn = received[15];			//Most significant bit is control bit
	 
	 //instantiate vga driver module
	 vga_core vga(clk,done,char,msgEn,clkdone,vgaclk,hsync,vsync,r,g,b);

endmodule

/////////////////////////////////////////////
// vga_spi
//   SPI slave interface is receive only
//   Instead of receiving a done bit, it just counts how many cycles of sck have occured
/////////////////////////////////////////////
module vga_spi(input logic sck, 		//From master
					input logic sdi,		//From master (is sdi)
					output logic done,	//done bit generated by counting
					output logic [15:0] q); // Data received
	
	//intermediate logic
	logic [6:0] counter;
	
	//spi shift register
	always_ff @(posedge sck)
		q <= {q[14:0], sdi}; 
	
	//done bit counter register
	always_ff@(posedge sck)
		if (counter == 16)
			counter <=1;
		else counter <= counter +1;
		
	//done when 16 bits have been received		
	assign done = (counter==16);
	
endmodule

///////////////////////////////////////////
// vga_core
// 	vga driver implementation
///////////////////////////////////////////
module vga_core(input logic clk,
					 input logic done,
					 input logic [7:0] char,
					 input logic msgEn,
					 output logic clkdone,
					 output logic vgaclk,
					 output logic hsync, vsync,
					 output logic r,g,b); //RGB values will be a single intensity
	//intermediate variables
	logic [9:0] x, y;		//x and ycounter
	logic [7:0] ch;		//character to be displayed
	
	// Using the wizard, PLL to create the 25.175 MHz VGA pixel clock
	// Screen is 800 clocks wide by 525 tall, but only 640 x 480 used
	// HSync = vgaclk/800 = 31.470 kHz
	// Vsync = Hsync / 525 = 59.94 Hz (~60 Hz refresh rate)
	//Hsync and Vsync dont have regular duty cycles, so have to do weird things
	PLLVGA PLLVGA_inst(.inclk0 ( clk ),.c0 ( vgaclk ));
		
	//instantiate character select module
	charSel msgShft(clk,done,clkdone,msgEn,char,x,y,ch);
	
	// Generate monitor timing signals
	vgaController vgaCont(vgaclk, hsync, vsync, x, y);
	
	// Module to determine whether pixels are on
	videoGen videoGen(x, y,ch, r, g, b);
	
endmodule

/////////////////////////////////////////////
// vgaController
//  vga implementation
/////////////////////////////////////////////
module vgaController #(parameter HBP = 10'd48,		  //H back porch
											HACTIVE = 10'd640,  //Horizontal active section
											HFP = 10'd16,		  //Horizontal front porch
											HSYN = 10'd96,		  //H sync time
											HMAX = HACTIVE + HFP + HSYN + HBP,
											VBP = 10'd32,
											VACTIVE = 10'd480,
											VFP = 10'd11,
											VSYN = 10'd2,
											VMAX = VACTIVE + VFP + VSYN + VBP)
							(input logic vgaclk,
							 output logic hsync, vsync, 
							 output logic [9:0] x, y); //10 bits for up to 1024 values
	// counters for horizontal and vertical positions
	always @(posedge vgaclk) begin
		x++;						//vga_clk iterates through pixels
		if (x == HMAX) begin	//If at last pixel, then we start over
			x = 0;
			y++;					//Increment row
			if (y == VMAX) 	//If last row, then start over
				y = 0;
			end
		end
	
	// Compute sync signals (active low (just not the output) Refer to pictures in Ch 9 of digital design
	assign hsync = ~(x >= HBP+ HACTIVE + HFP & x < HMAX);
	assign vsync = ~(y >= VBP+ VACTIVE + VFP & y < VMAX);

endmodule

/////////////////////////////////////////////
// videogen
//  vga implementation
/////////////////////////////////////////////
module videoGen(input logic [9:0] x, y, 
					 input logic [7:0] ch, 
					 output logic r,g,b);
	logic pixelOn;
	// Given y position, choose a character to display
	// then look up the pixel value from the character ROM
	// and display it in red or blue.Also draw a green rectangle.
	chargenrom charrom_inst(ch, x[5:0], y[5:0], pixelOn);
	
	assign r =pixelOn;
	assign g =pixelOn;
	assign b =pixelOn;
	
endmodule

/////////////////////////////////////////////
// chargenrom
//  vga implementation
/////////////////////////////////////////////
module chargenrom(input logic [7:0] ch, //ascii value
						input logic [5:0] xoff, yoff,
						output logic pixelOn);
	logic [31:0] charrom[26623:0]; // character generator ROM only need 6 bits
	logic [31:0] line; // a line read from the ROM
	
	// Initialize ROM with characters from text file
	initial
		$readmemb("char.txt", charrom);
	
	// Index into ROM to find line of character
	assign line = charrom[yoff + {ch-65,5'b00000}]; // Subtract 65 because A
																  // is entry 0
	// Reverse order of bits when picking
	//Left most col in ROM is most significant
	//Drawn in least significant x position
	assign pixelOn = line[5'd31-xoff];
	
endmodule

module megaflop(input logic clk,
					 input logic done,
					 input logic en,
					 input logic [7:0] ch,
					 output logic [7:0] q0,q1,q2,q3,q4,q5,q6,q7,q8,q9,q10,q11,q12,q13,q14 );
	 always_ff@(posedge clk)
		if(done&en) 
			begin
					q0 <= ch;
					q1 <= q0;
					q2 <= q1;
					q3 <= q2;
					q4 <= q3;
					q5 <= q4;
					q6 <= q5;
					q7 <= q6;
					q8 <= q7;
					q9 <= q8;
					q10<= q9;
					q11 <= q10;
					q12 <= q11;
					q13 <= q12;
					q14 <= q13;
			end
endmodule

module charSel #(parameter CHW = 10'd32,
								  CHH = 10'd32,
								  HBP = 10'd48,		  //H back porch
								  HACTIVE = 10'd640,  //Horizontal active section
								  HFP = 10'd16,		  //Horizontal front porch
								  HSYN = 10'd96,		  //H sync time
								  HMAX = HACTIVE + HFP + HSYN + HBP,
								  VBP = 10'd32,
								  VACTIVE = 10'd480,
								  VFP = 10'd11,
								  VSYN = 10'd2,
								  VMAX = VACTIVE + VFP + VSYN + VBP)
				 (input logic clk,
				  input logic done,
				  output logic clkdone,
				  input logic msgEn,
				  input logic [7:0] char,
				  input logic [9:0] x,y,
				  output logic [7:0] ch);
	  
	  logic [7:0] m0,m1,m2,m3,m4,m5,m6,m7,m8,m9,m10,m11,m12,m13,m14;
	  logic [7:0] l0,l1,l2,l3,l4,l5,l6,l7,l8,l9,l10,l11,l12,l13,l14;
	  logic hasntdone; 
	  always_ff@(posedge clk)
	   if (~done) 
			begin 
			clkdone<=0;
			hasntdone<=1;
			end
		else if (hasntdone&done) 
		begin
			hasntdone<=0;
			clkdone<=1;
		end
		else clkdone<=0;
			
	  megaflop msg_flop(clk,clkdone,msgEn,char,m0,m1,m2,m3,m4,m5,m6,m7,m8,m9,m10,m11,m12,m13,m14);
	  
	  
	  megaflop loc_flop(clk,clkdone,~msgEn,char,l0,l1,l2,l3,l4,l5,l6,l7,l8,l9,l10,l11,l12,l13,l14);
	  

	  logic[7:0] chm,chl;
	  charLocX locxm(x,m0,m1,m2,m3,m4,m5,m6,m7,m8,m9,m10,m11,m12,m13,m14,chm);
	  
	  charLocX locxl(x,l0,l1,l2,l3,l4,l5,l6,l7,l8,l9,l10,l11,l12,l13,l14,chl);
	  charLocY locy(y,chm,chl,ch);
	  		
endmodule

module charLocX #(parameter CHW = 10'd32,
								  CHH = 10'd32,
								  HBP = 10'd48,		  //H back porch
								  HACTIVE = 10'd640,  //Horizontal active section
								  HFP = 10'd16,		  //Horizontal front porch
								  HSYN = 10'd96,		  //H sync time
								  HMAX = HACTIVE + HFP + HSYN + HBP,
								  VBP = 10'd32,
								  VACTIVE = 10'd480,
								  VFP = 10'd11,
								  VSYN = 10'd2,
								  VMAX = VACTIVE + VFP + VSYN + VBP)
				 
				 (input logic [9:0] x,
				  input logic [7:0] m0,m1,m2,m3,m4,m5,m6,m7,m8,m9,m10,m11,m12,m13,m14,
				  output logic [7:0] ch);
				  
	  always_comb
		if		 (0<x&x<3*CHW ) 		  ch=00;
		else if((4*CHW<x) & (x<(5*CHW-1))) ch=m0; //Dont do <= this gets rid of overlap
		else if((5*CHW<x) & (x<(6*CHW-1))) ch=m1;
		else if((6*CHW<x) & (x<(7*CHW-1))) ch=m2;
		else if((7*CHW<x) & (x<(8*CHW-1))) ch=m3;
		else if((8*CHW<x) & (x<(9*CHW-1))) ch=m4;
		else if((9*CHW<x) & (x<(10*CHW-1))) ch=m5;
		else if((10*CHW<x) & (x<(11*CHW-1))) ch=m6;
		else if((11*CHW<x) & (x<(12*CHW-1))) ch=m7;
		else if((12*CHW<x) & (x<(13*CHW-1))) ch=m8;
		else if((13*CHW<x) & (x<(14*CHW-1))) ch=m9;
		else if((14*CHW<x) & (x<(15*CHW-1))) ch=m10;
		else if((15*CHW<x) & (x<(16*CHW-1))) ch=m11;
		else if((16*CHW<x) & (x<(17*CHW-1))) ch=m12;
		else if((17*CHW<x) & (x<(18*CHW-1))) ch=m13;
		else if((18*CHW<x) & (x<(19*CHW-1))) ch=m14;
		else ch=00;		
endmodule	

module charLocY #(parameter CHW = 10'd32,
								  CHH = 10'd32,
								  HBP = 10'd48,		  //H back porch
								  HACTIVE = 10'd640,  //Horizontal active section
								  HFP = 10'd16,		  //Horizontal front porch
								  HSYN = 10'd96,		  //H sync time
								  HMAX = HACTIVE + HFP + HSYN + HBP,
								  VBP = 10'd32,
								  VACTIVE = 10'd480,
								  VFP = 10'd11,
								  VSYN = 10'd2,
								  VMAX = VACTIVE + VFP + VSYN + VBP)
				 (input logic [9:0] y,
				  input logic [7:0] chm, chl,
				  output logic [7:0] ch);
				  
	  always_comb
		if		 (0<y&y<3*CHH ) 		  ch=00;
		else if((4*CHH<=y) & (y<(5*CHH))) ch=chm;
		else if((8*CHH<=y) & (y<(9*CHH))) ch=chl;
		else ch=00;		
endmodule
  

